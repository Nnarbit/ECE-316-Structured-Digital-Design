library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.numeric_std.all;

entity ALUB is
	port (Din : in std_logic_vector(9 downto 0); 
		LoadX, LoadY, Clk : in std_logic;
		Dout0, Dout1 : out std_logic_vector(6 downto 0);
		Overflow, Negative: out std_logic);
end ALUB;

architecture struct of ALUB is
   component reg8 is
	Port(Clk : in std_logic;
           Input : in  std_logic_vector (7 downto 0);
           Load : in  std_logic;
           Output : out  std_logic_vector (7 downto 0));
   end component;

   component addo is
	   port (A, B : in  std_logic_vector(7 downto 0);
		Opr : in std_logic_vector(2 downto 0);
		Dout : out std_logic_vector(7 downto 0);
		Overflow, Negative: out std_logic);
   end component;

   component BCD is
	   port (Din: in std_logic_vector(7 downto 0);
		 D0out, D1out: out std_logic_vector(3 downto 0);
	         overflow: out std_logic);
   end component;
	
   component sevensegdisplay is 
	   port(A, B, C, D : in std_logic;
      		Sa, Sb, Sc, Sd, Se, Sf, Sg : out std_logic);
   end component;

  Signal Rx : std_logic_vector(7 downto 0);
  Signal Ry : std_logic_vector(7 downto 0);
  Signal Sum : std_logic_vector(7 downto 0);	
  Signal Bx : std_logic_vector(3 downto 0);
  Signal By: std_logic_vector(3 downto 0);
  Signal OvF: std_logic;

begin
  RegX: reg8 port map(Clk, Din(7 downto 0), LoadX, Rx);
  RegY: reg8 port map(Clk, Din(7 downto 0), LoadY, Ry);
  Adder: addo port map(Rx, Ry, Din(9 downto 7), Sum, Overflow, Negative);
  B_C_D: BCD port map(Sum, Bx, By, OvF);
  dispx: sevensegdisplay port map(Bx(3), Bx(2), Bx(1), Bx(0), Dout0(0), Dout0(1), Dout0(2), Dout0(3), Dout0(4), Dout0(5), Dout0(6));
  dispy: sevensegdisplay port map(By(3), By(2), By(1), By(0), Dout1(0), Dout1(1), Dout1(2), Dout1(3), Dout1(4), Dout1(5), Dout1(6));
  
end struct;
